/*
    Created             : /home/caonam/SNN_THESIS_PROJECT/RTL/ADDER.v
    Module Name         : ADDER
    Author              : Van Nam CAO
    Date                : 08 - 07 - 2025
    Description         : This module that perform 32-bit floating point addition
*/

module ADDER (
    // FIXME: define ports
);

endmodule
